`ifndef DESINES_SVH_
`define DESINES_SVH_

`include "scr1_arch_description.svh"
`include "scr1_arch_types.svh"

`define LANE 16
 typedef  type_scr1_mprf_v[`LANE - 1 : 0] type_vector;



`endif
